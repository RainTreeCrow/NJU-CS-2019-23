module level_text_setter(clk, game_reset, inlevelDisplay, current_level, main_difficulty, x_pointer, y_pointer, level_text, finished_displaying_level);
// display for 3 seconds!
	input game_reset;
   input inlevelDisplay;
	input [3:0] main_difficulty;
	input [3:0] current_level;
   input clk;
   input [7:0]x_pointer;
	input [6:0]y_pointer;
	output reg level_text; // check if the pixel is the menu's text.
	output reg finished_displaying_level;
	
	reg [31:0] counter;
	
	//countdown
	always@(posedge clk)
	begin
		if (game_reset)
			counter = 149999999;
		if (inlevelDisplay) begin
			if (counter == 0)
				counter = 149999999;
			counter = counter - 1;
		finished_displaying_level = counter == 0 ? 1 : 0;
		end
	end
	

	//menu's normal text
	always@(posedge clk)
	begin
		if (inlevelDisplay)
			 begin
			 if (main_texts || difficulty_display || level_display)
				 level_text <= 1'b1;
			 else
				 level_text <= 1'b0;
			 end
	end

	wire main_texts = (x_pointer == 54 && y_pointer == 41)
||(x_pointer == 55 && y_pointer == 41)
||(x_pointer == 61 && y_pointer == 41)
||(x_pointer == 62 && y_pointer == 41)
||(x_pointer == 63 && y_pointer == 41)
||(x_pointer == 64 && y_pointer == 41)
||(x_pointer == 65 && y_pointer == 41)
||(x_pointer == 66 && y_pointer == 41)
||(x_pointer == 68 && y_pointer == 41)
||(x_pointer == 69 && y_pointer == 41)
||(x_pointer == 73 && y_pointer == 41)
||(x_pointer == 74 && y_pointer == 41)
||(x_pointer == 76 && y_pointer == 41)
||(x_pointer == 77 && y_pointer == 41)
||(x_pointer == 78 && y_pointer == 41)
||(x_pointer == 79 && y_pointer == 41)
||(x_pointer == 80 && y_pointer == 41)
||(x_pointer == 81 && y_pointer == 41)
||(x_pointer == 83 && y_pointer == 41)
||(x_pointer == 84 && y_pointer == 41)
||(x_pointer == 54 && y_pointer == 42)
||(x_pointer == 55 && y_pointer == 42)
||(x_pointer == 61 && y_pointer == 42)
||(x_pointer == 62 && y_pointer == 42)
||(x_pointer == 68 && y_pointer == 42)
||(x_pointer == 69 && y_pointer == 42)
||(x_pointer == 73 && y_pointer == 42)
||(x_pointer == 74 && y_pointer == 42)
||(x_pointer == 76 && y_pointer == 42)
||(x_pointer == 77 && y_pointer == 42)
||(x_pointer == 83 && y_pointer == 42)
||(x_pointer == 84 && y_pointer == 42)
||(x_pointer == 54 && y_pointer == 43)
||(x_pointer == 55 && y_pointer == 43)
||(x_pointer == 61 && y_pointer == 43)
||(x_pointer == 62 && y_pointer == 43)
||(x_pointer == 68 && y_pointer == 43)
||(x_pointer == 69 && y_pointer == 43)
||(x_pointer == 73 && y_pointer == 43)
||(x_pointer == 74 && y_pointer == 43)
||(x_pointer == 76 && y_pointer == 43)
||(x_pointer == 77 && y_pointer == 43)
||(x_pointer == 83 && y_pointer == 43)
||(x_pointer == 84 && y_pointer == 43)
||(x_pointer == 54 && y_pointer == 44)
||(x_pointer == 55 && y_pointer == 44)
||(x_pointer == 61 && y_pointer == 44)
||(x_pointer == 62 && y_pointer == 44)
||(x_pointer == 69 && y_pointer == 44)
||(x_pointer == 70 && y_pointer == 44)
||(x_pointer == 72 && y_pointer == 44)
||(x_pointer == 73 && y_pointer == 44)
||(x_pointer == 74 && y_pointer == 44)
||(x_pointer == 76 && y_pointer == 44)
||(x_pointer == 77 && y_pointer == 44)
||(x_pointer == 83 && y_pointer == 44)
||(x_pointer == 84 && y_pointer == 44)
||(x_pointer == 54 && y_pointer == 45)
||(x_pointer == 55 && y_pointer == 45)
||(x_pointer == 61 && y_pointer == 45)
||(x_pointer == 62 && y_pointer == 45)
||(x_pointer == 69 && y_pointer == 45)
||(x_pointer == 70 && y_pointer == 45)
||(x_pointer == 72 && y_pointer == 45)
||(x_pointer == 73 && y_pointer == 45)
||(x_pointer == 76 && y_pointer == 45)
||(x_pointer == 77 && y_pointer == 45)
||(x_pointer == 83 && y_pointer == 45)
||(x_pointer == 84 && y_pointer == 45)
||(x_pointer == 54 && y_pointer == 46)
||(x_pointer == 55 && y_pointer == 46)
||(x_pointer == 61 && y_pointer == 46)
||(x_pointer == 62 && y_pointer == 46)
||(x_pointer == 63 && y_pointer == 46)
||(x_pointer == 64 && y_pointer == 46)
||(x_pointer == 65 && y_pointer == 46)
||(x_pointer == 66 && y_pointer == 46)
||(x_pointer == 69 && y_pointer == 46)
||(x_pointer == 70 && y_pointer == 46)
||(x_pointer == 71 && y_pointer == 46)
||(x_pointer == 72 && y_pointer == 46)
||(x_pointer == 73 && y_pointer == 46)
||(x_pointer == 76 && y_pointer == 46)
||(x_pointer == 77 && y_pointer == 46)
||(x_pointer == 78 && y_pointer == 46)
||(x_pointer == 79 && y_pointer == 46)
||(x_pointer == 80 && y_pointer == 46)
||(x_pointer == 81 && y_pointer == 46)
||(x_pointer == 83 && y_pointer == 46)
||(x_pointer == 84 && y_pointer == 46)
||(x_pointer == 54 && y_pointer == 47)
||(x_pointer == 55 && y_pointer == 47)
||(x_pointer == 61 && y_pointer == 47)
||(x_pointer == 62 && y_pointer == 47)
||(x_pointer == 69 && y_pointer == 47)
||(x_pointer == 70 && y_pointer == 47)
||(x_pointer == 71 && y_pointer == 47)
||(x_pointer == 72 && y_pointer == 47)
||(x_pointer == 73 && y_pointer == 47)
||(x_pointer == 76 && y_pointer == 47)
||(x_pointer == 77 && y_pointer == 47)
||(x_pointer == 83 && y_pointer == 47)
||(x_pointer == 84 && y_pointer == 47)
||(x_pointer == 54 && y_pointer == 48)
||(x_pointer == 55 && y_pointer == 48)
||(x_pointer == 61 && y_pointer == 48)
||(x_pointer == 62 && y_pointer == 48)
||(x_pointer == 70 && y_pointer == 48)
||(x_pointer == 71 && y_pointer == 48)
||(x_pointer == 72 && y_pointer == 48)
||(x_pointer == 76 && y_pointer == 48)
||(x_pointer == 77 && y_pointer == 48)
||(x_pointer == 83 && y_pointer == 48)
||(x_pointer == 84 && y_pointer == 48)
||(x_pointer == 54 && y_pointer == 49)
||(x_pointer == 55 && y_pointer == 49)
||(x_pointer == 61 && y_pointer == 49)
||(x_pointer == 62 && y_pointer == 49)
||(x_pointer == 70 && y_pointer == 49)
||(x_pointer == 71 && y_pointer == 49)
||(x_pointer == 72 && y_pointer == 49)
||(x_pointer == 76 && y_pointer == 49)
||(x_pointer == 77 && y_pointer == 49)
||(x_pointer == 83 && y_pointer == 49)
||(x_pointer == 84 && y_pointer == 49)
||(x_pointer == 54 && y_pointer == 50)
||(x_pointer == 55 && y_pointer == 50)
||(x_pointer == 61 && y_pointer == 50)
||(x_pointer == 62 && y_pointer == 50)
||(x_pointer == 71 && y_pointer == 50)
||(x_pointer == 76 && y_pointer == 50)
||(x_pointer == 77 && y_pointer == 50)
||(x_pointer == 83 && y_pointer == 50)
||(x_pointer == 84 && y_pointer == 50)
||(x_pointer == 54 && y_pointer == 51)
||(x_pointer == 55 && y_pointer == 51)
||(x_pointer == 56 && y_pointer == 51)
||(x_pointer == 57 && y_pointer == 51)
||(x_pointer == 58 && y_pointer == 51)
||(x_pointer == 59 && y_pointer == 51)
||(x_pointer == 61 && y_pointer == 51)
||(x_pointer == 62 && y_pointer == 51)
||(x_pointer == 63 && y_pointer == 51)
||(x_pointer == 64 && y_pointer == 51)
||(x_pointer == 65 && y_pointer == 51)
||(x_pointer == 66 && y_pointer == 51)
||(x_pointer == 71 && y_pointer == 51)
||(x_pointer == 76 && y_pointer == 51)
||(x_pointer == 77 && y_pointer == 51)
||(x_pointer == 78 && y_pointer == 51)
||(x_pointer == 79 && y_pointer == 51)
||(x_pointer == 80 && y_pointer == 51)
||(x_pointer == 81 && y_pointer == 51)
||(x_pointer == 83 && y_pointer == 51)
||(x_pointer == 84 && y_pointer == 51)
||(x_pointer == 85 && y_pointer == 51)
||(x_pointer == 86 && y_pointer == 51)
||(x_pointer == 87 && y_pointer == 51)
||(x_pointer == 88 && y_pointer == 51);


	wire difficulty_display = (main_difficulty == 4'd4 && ((x_pointer == 62 && y_pointer == 65)
||(x_pointer == 63 && y_pointer == 65)
||(x_pointer == 64 && y_pointer == 65)
||(x_pointer == 65 && y_pointer == 65)
||(x_pointer == 66 && y_pointer == 65)
||(x_pointer == 67 && y_pointer == 65)
||(x_pointer == 71 && y_pointer == 65)
||(x_pointer == 72 && y_pointer == 65)
||(x_pointer == 73 && y_pointer == 65)
||(x_pointer == 78 && y_pointer == 65)
||(x_pointer == 79 && y_pointer == 65)
||(x_pointer == 80 && y_pointer == 65)
||(x_pointer == 81 && y_pointer == 65)
||(x_pointer == 82 && y_pointer == 65)
||(x_pointer == 83 && y_pointer == 65)
||(x_pointer == 85 && y_pointer == 65)
||(x_pointer == 86 && y_pointer == 65)
||(x_pointer == 91 && y_pointer == 65)
||(x_pointer == 92 && y_pointer == 65)
||(x_pointer == 62 && y_pointer == 66)
||(x_pointer == 63 && y_pointer == 66)
||(x_pointer == 71 && y_pointer == 66)
||(x_pointer == 72 && y_pointer == 66)
||(x_pointer == 73 && y_pointer == 66)
||(x_pointer == 77 && y_pointer == 66)
||(x_pointer == 78 && y_pointer == 66)
||(x_pointer == 82 && y_pointer == 66)
||(x_pointer == 83 && y_pointer == 66)
||(x_pointer == 85 && y_pointer == 66)
||(x_pointer == 86 && y_pointer == 66)
||(x_pointer == 91 && y_pointer == 66)
||(x_pointer == 92 && y_pointer == 66)
||(x_pointer == 62 && y_pointer == 67)
||(x_pointer == 63 && y_pointer == 67)
||(x_pointer == 71 && y_pointer == 67)
||(x_pointer == 72 && y_pointer == 67)
||(x_pointer == 73 && y_pointer == 67)
||(x_pointer == 77 && y_pointer == 67)
||(x_pointer == 78 && y_pointer == 67)
||(x_pointer == 82 && y_pointer == 67)
||(x_pointer == 83 && y_pointer == 67)
||(x_pointer == 86 && y_pointer == 67)
||(x_pointer == 87 && y_pointer == 67)
||(x_pointer == 90 && y_pointer == 67)
||(x_pointer == 91 && y_pointer == 67)
||(x_pointer == 62 && y_pointer == 68)
||(x_pointer == 63 && y_pointer == 68)
||(x_pointer == 71 && y_pointer == 68)
||(x_pointer == 73 && y_pointer == 68)
||(x_pointer == 77 && y_pointer == 68)
||(x_pointer == 78 && y_pointer == 68)
||(x_pointer == 79 && y_pointer == 68)
||(x_pointer == 82 && y_pointer == 68)
||(x_pointer == 83 && y_pointer == 68)
||(x_pointer == 86 && y_pointer == 68)
||(x_pointer == 87 && y_pointer == 68)
||(x_pointer == 88 && y_pointer == 68)
||(x_pointer == 89 && y_pointer == 68)
||(x_pointer == 90 && y_pointer == 68)
||(x_pointer == 91 && y_pointer == 68)
||(x_pointer == 62 && y_pointer == 69)
||(x_pointer == 63 && y_pointer == 69)
||(x_pointer == 71 && y_pointer == 69)
||(x_pointer == 73 && y_pointer == 69)
||(x_pointer == 78 && y_pointer == 69)
||(x_pointer == 79 && y_pointer == 69)
||(x_pointer == 80 && y_pointer == 69)
||(x_pointer == 87 && y_pointer == 69)
||(x_pointer == 88 && y_pointer == 69)
||(x_pointer == 89 && y_pointer == 69)
||(x_pointer == 90 && y_pointer == 69)
||(x_pointer == 62 && y_pointer == 70)
||(x_pointer == 63 && y_pointer == 70)
||(x_pointer == 64 && y_pointer == 70)
||(x_pointer == 65 && y_pointer == 70)
||(x_pointer == 66 && y_pointer == 70)
||(x_pointer == 67 && y_pointer == 70)
||(x_pointer == 70 && y_pointer == 70)
||(x_pointer == 71 && y_pointer == 70)
||(x_pointer == 73 && y_pointer == 70)
||(x_pointer == 74 && y_pointer == 70)
||(x_pointer == 79 && y_pointer == 70)
||(x_pointer == 80 && y_pointer == 70)
||(x_pointer == 81 && y_pointer == 70)
||(x_pointer == 87 && y_pointer == 70)
||(x_pointer == 88 && y_pointer == 70)
||(x_pointer == 89 && y_pointer == 70)
||(x_pointer == 90 && y_pointer == 70)
||(x_pointer == 62 && y_pointer == 71)
||(x_pointer == 63 && y_pointer == 71)
||(x_pointer == 70 && y_pointer == 71)
||(x_pointer == 71 && y_pointer == 71)
||(x_pointer == 73 && y_pointer == 71)
||(x_pointer == 74 && y_pointer == 71)
||(x_pointer == 80 && y_pointer == 71)
||(x_pointer == 81 && y_pointer == 71)
||(x_pointer == 82 && y_pointer == 71)
||(x_pointer == 88 && y_pointer == 71)
||(x_pointer == 89 && y_pointer == 71)
||(x_pointer == 62 && y_pointer == 72)
||(x_pointer == 63 && y_pointer == 72)
||(x_pointer == 70 && y_pointer == 72)
||(x_pointer == 71 && y_pointer == 72)
||(x_pointer == 72 && y_pointer == 72)
||(x_pointer == 73 && y_pointer == 72)
||(x_pointer == 74 && y_pointer == 72)
||(x_pointer == 81 && y_pointer == 72)
||(x_pointer == 82 && y_pointer == 72)
||(x_pointer == 83 && y_pointer == 72)
||(x_pointer == 88 && y_pointer == 72)
||(x_pointer == 89 && y_pointer == 72)
||(x_pointer == 62 && y_pointer == 73)
||(x_pointer == 63 && y_pointer == 73)
||(x_pointer == 70 && y_pointer == 73)
||(x_pointer == 71 && y_pointer == 73)
||(x_pointer == 72 && y_pointer == 73)
||(x_pointer == 73 && y_pointer == 73)
||(x_pointer == 74 && y_pointer == 73)
||(x_pointer == 82 && y_pointer == 73)
||(x_pointer == 83 && y_pointer == 73)
||(x_pointer == 88 && y_pointer == 73)
||(x_pointer == 89 && y_pointer == 73)
||(x_pointer == 62 && y_pointer == 74)
||(x_pointer == 63 && y_pointer == 74)
||(x_pointer == 69 && y_pointer == 74)
||(x_pointer == 70 && y_pointer == 74)
||(x_pointer == 74 && y_pointer == 74)
||(x_pointer == 75 && y_pointer == 74)
||(x_pointer == 77 && y_pointer == 74)
||(x_pointer == 78 && y_pointer == 74)
||(x_pointer == 82 && y_pointer == 74)
||(x_pointer == 83 && y_pointer == 74)
||(x_pointer == 88 && y_pointer == 74)
||(x_pointer == 89 && y_pointer == 74)
||(x_pointer == 62 && y_pointer == 75)
||(x_pointer == 63 && y_pointer == 75)
||(x_pointer == 69 && y_pointer == 75)
||(x_pointer == 70 && y_pointer == 75)
||(x_pointer == 74 && y_pointer == 75)
||(x_pointer == 75 && y_pointer == 75)
||(x_pointer == 77 && y_pointer == 75)
||(x_pointer == 78 && y_pointer == 75)
||(x_pointer == 82 && y_pointer == 75)
||(x_pointer == 83 && y_pointer == 75)
||(x_pointer == 88 && y_pointer == 75)
||(x_pointer == 89 && y_pointer == 75)
||(x_pointer == 62 && y_pointer == 76)
||(x_pointer == 63 && y_pointer == 76)
||(x_pointer == 64 && y_pointer == 76)
||(x_pointer == 65 && y_pointer == 76)
||(x_pointer == 66 && y_pointer == 76)
||(x_pointer == 67 && y_pointer == 76)
||(x_pointer == 69 && y_pointer == 76)
||(x_pointer == 70 && y_pointer == 76)
||(x_pointer == 74 && y_pointer == 76)
||(x_pointer == 75 && y_pointer == 76)
||(x_pointer == 78 && y_pointer == 76)
||(x_pointer == 79 && y_pointer == 76)
||(x_pointer == 80 && y_pointer == 76)
||(x_pointer == 81 && y_pointer == 76)
||(x_pointer == 82 && y_pointer == 76)
||(x_pointer == 83 && y_pointer == 76)
||(x_pointer == 88 && y_pointer == 76)
||(x_pointer == 89 && y_pointer == 76))) || (main_difficulty == 4'd2 && ((x_pointer == 54 && y_pointer == 65)
||(x_pointer == 55 && y_pointer == 65)
||(x_pointer == 59 && y_pointer == 65)
||(x_pointer == 60 && y_pointer == 65)
||(x_pointer == 62 && y_pointer == 65)
||(x_pointer == 63 && y_pointer == 65)
||(x_pointer == 64 && y_pointer == 65)
||(x_pointer == 65 && y_pointer == 65)
||(x_pointer == 66 && y_pointer == 65)
||(x_pointer == 67 && y_pointer == 65)
||(x_pointer == 68 && y_pointer == 65)
||(x_pointer == 69 && y_pointer == 65)
||(x_pointer == 71 && y_pointer == 65)
||(x_pointer == 72 && y_pointer == 65)
||(x_pointer == 73 && y_pointer == 65)
||(x_pointer == 74 && y_pointer == 65)
||(x_pointer == 75 && y_pointer == 65)
||(x_pointer == 76 && y_pointer == 65)
||(x_pointer == 77 && y_pointer == 65)
||(x_pointer == 80 && y_pointer == 65)
||(x_pointer == 81 && y_pointer == 65)
||(x_pointer == 86 && y_pointer == 65)
||(x_pointer == 87 && y_pointer == 65)
||(x_pointer == 91 && y_pointer == 65)
||(x_pointer == 92 && y_pointer == 65)
||(x_pointer == 93 && y_pointer == 65)
||(x_pointer == 97 && y_pointer == 65)
||(x_pointer == 98 && y_pointer == 65)
||(x_pointer == 54 && y_pointer == 66)
||(x_pointer == 55 && y_pointer == 66)
||(x_pointer == 59 && y_pointer == 66)
||(x_pointer == 60 && y_pointer == 66)
||(x_pointer == 62 && y_pointer == 66)
||(x_pointer == 63 && y_pointer == 66)
||(x_pointer == 68 && y_pointer == 66)
||(x_pointer == 69 && y_pointer == 66)
||(x_pointer == 71 && y_pointer == 66)
||(x_pointer == 72 && y_pointer == 66)
||(x_pointer == 76 && y_pointer == 66)
||(x_pointer == 77 && y_pointer == 66)
||(x_pointer == 80 && y_pointer == 66)
||(x_pointer == 81 && y_pointer == 66)
||(x_pointer == 86 && y_pointer == 66)
||(x_pointer == 87 && y_pointer == 66)
||(x_pointer == 91 && y_pointer == 66)
||(x_pointer == 92 && y_pointer == 66)
||(x_pointer == 93 && y_pointer == 66)
||(x_pointer == 97 && y_pointer == 66)
||(x_pointer == 98 && y_pointer == 66)
||(x_pointer == 54 && y_pointer == 67)
||(x_pointer == 55 && y_pointer == 67)
||(x_pointer == 59 && y_pointer == 67)
||(x_pointer == 60 && y_pointer == 67)
||(x_pointer == 62 && y_pointer == 67)
||(x_pointer == 63 && y_pointer == 67)
||(x_pointer == 68 && y_pointer == 67)
||(x_pointer == 69 && y_pointer == 67)
||(x_pointer == 71 && y_pointer == 67)
||(x_pointer == 72 && y_pointer == 67)
||(x_pointer == 76 && y_pointer == 67)
||(x_pointer == 77 && y_pointer == 67)
||(x_pointer == 80 && y_pointer == 67)
||(x_pointer == 81 && y_pointer == 67)
||(x_pointer == 82 && y_pointer == 67)
||(x_pointer == 85 && y_pointer == 67)
||(x_pointer == 86 && y_pointer == 67)
||(x_pointer == 87 && y_pointer == 67)
||(x_pointer == 91 && y_pointer == 67)
||(x_pointer == 92 && y_pointer == 67)
||(x_pointer == 93 && y_pointer == 67)
||(x_pointer == 97 && y_pointer == 67)
||(x_pointer == 98 && y_pointer == 67)
||(x_pointer == 54 && y_pointer == 68)
||(x_pointer == 55 && y_pointer == 68)
||(x_pointer == 56 && y_pointer == 68)
||(x_pointer == 59 && y_pointer == 68)
||(x_pointer == 60 && y_pointer == 68)
||(x_pointer == 62 && y_pointer == 68)
||(x_pointer == 63 && y_pointer == 68)
||(x_pointer == 68 && y_pointer == 68)
||(x_pointer == 69 && y_pointer == 68)
||(x_pointer == 71 && y_pointer == 68)
||(x_pointer == 72 && y_pointer == 68)
||(x_pointer == 76 && y_pointer == 68)
||(x_pointer == 77 && y_pointer == 68)
||(x_pointer == 80 && y_pointer == 68)
||(x_pointer == 81 && y_pointer == 68)
||(x_pointer == 82 && y_pointer == 68)
||(x_pointer == 85 && y_pointer == 68)
||(x_pointer == 86 && y_pointer == 68)
||(x_pointer == 87 && y_pointer == 68)
||(x_pointer == 91 && y_pointer == 68)
||(x_pointer == 93 && y_pointer == 68)
||(x_pointer == 97 && y_pointer == 68)
||(x_pointer == 98 && y_pointer == 68)
||(x_pointer == 54 && y_pointer == 69)
||(x_pointer == 55 && y_pointer == 69)
||(x_pointer == 56 && y_pointer == 69)
||(x_pointer == 59 && y_pointer == 69)
||(x_pointer == 60 && y_pointer == 69)
||(x_pointer == 62 && y_pointer == 69)
||(x_pointer == 63 && y_pointer == 69)
||(x_pointer == 68 && y_pointer == 69)
||(x_pointer == 69 && y_pointer == 69)
||(x_pointer == 71 && y_pointer == 69)
||(x_pointer == 72 && y_pointer == 69)
||(x_pointer == 76 && y_pointer == 69)
||(x_pointer == 77 && y_pointer == 69)
||(x_pointer == 80 && y_pointer == 69)
||(x_pointer == 81 && y_pointer == 69)
||(x_pointer == 82 && y_pointer == 69)
||(x_pointer == 85 && y_pointer == 69)
||(x_pointer == 86 && y_pointer == 69)
||(x_pointer == 87 && y_pointer == 69)
||(x_pointer == 91 && y_pointer == 69)
||(x_pointer == 93 && y_pointer == 69)
||(x_pointer == 97 && y_pointer == 69)
||(x_pointer == 98 && y_pointer == 69)
||(x_pointer == 54 && y_pointer == 70)
||(x_pointer == 55 && y_pointer == 70)
||(x_pointer == 56 && y_pointer == 70)
||(x_pointer == 57 && y_pointer == 70)
||(x_pointer == 59 && y_pointer == 70)
||(x_pointer == 60 && y_pointer == 70)
||(x_pointer == 62 && y_pointer == 70)
||(x_pointer == 63 && y_pointer == 70)
||(x_pointer == 68 && y_pointer == 70)
||(x_pointer == 69 && y_pointer == 70)
||(x_pointer == 71 && y_pointer == 70)
||(x_pointer == 72 && y_pointer == 70)
||(x_pointer == 73 && y_pointer == 70)
||(x_pointer == 74 && y_pointer == 70)
||(x_pointer == 75 && y_pointer == 70)
||(x_pointer == 76 && y_pointer == 70)
||(x_pointer == 77 && y_pointer == 70)
||(x_pointer == 80 && y_pointer == 70)
||(x_pointer == 81 && y_pointer == 70)
||(x_pointer == 82 && y_pointer == 70)
||(x_pointer == 85 && y_pointer == 70)
||(x_pointer == 86 && y_pointer == 70)
||(x_pointer == 87 && y_pointer == 70)
||(x_pointer == 90 && y_pointer == 70)
||(x_pointer == 91 && y_pointer == 70)
||(x_pointer == 93 && y_pointer == 70)
||(x_pointer == 94 && y_pointer == 70)
||(x_pointer == 97 && y_pointer == 70)
||(x_pointer == 98 && y_pointer == 70)
||(x_pointer == 54 && y_pointer == 71)
||(x_pointer == 55 && y_pointer == 71)
||(x_pointer == 56 && y_pointer == 71)
||(x_pointer == 57 && y_pointer == 71)
||(x_pointer == 59 && y_pointer == 71)
||(x_pointer == 60 && y_pointer == 71)
||(x_pointer == 62 && y_pointer == 71)
||(x_pointer == 63 && y_pointer == 71)
||(x_pointer == 68 && y_pointer == 71)
||(x_pointer == 69 && y_pointer == 71)
||(x_pointer == 71 && y_pointer == 71)
||(x_pointer == 72 && y_pointer == 71)
||(x_pointer == 74 && y_pointer == 71)
||(x_pointer == 75 && y_pointer == 71)
||(x_pointer == 80 && y_pointer == 71)
||(x_pointer == 81 && y_pointer == 71)
||(x_pointer == 82 && y_pointer == 71)
||(x_pointer == 83 && y_pointer == 71)
||(x_pointer == 84 && y_pointer == 71)
||(x_pointer == 85 && y_pointer == 71)
||(x_pointer == 86 && y_pointer == 71)
||(x_pointer == 87 && y_pointer == 71)
||(x_pointer == 90 && y_pointer == 71)
||(x_pointer == 91 && y_pointer == 71)
||(x_pointer == 93 && y_pointer == 71)
||(x_pointer == 94 && y_pointer == 71)
||(x_pointer == 97 && y_pointer == 71)
||(x_pointer == 98 && y_pointer == 71)
||(x_pointer == 54 && y_pointer == 72)
||(x_pointer == 55 && y_pointer == 72)
||(x_pointer == 57 && y_pointer == 72)
||(x_pointer == 58 && y_pointer == 72)
||(x_pointer == 59 && y_pointer == 72)
||(x_pointer == 60 && y_pointer == 72)
||(x_pointer == 62 && y_pointer == 72)
||(x_pointer == 63 && y_pointer == 72)
||(x_pointer == 68 && y_pointer == 72)
||(x_pointer == 69 && y_pointer == 72)
||(x_pointer == 71 && y_pointer == 72)
||(x_pointer == 72 && y_pointer == 72)
||(x_pointer == 74 && y_pointer == 72)
||(x_pointer == 75 && y_pointer == 72)
||(x_pointer == 80 && y_pointer == 72)
||(x_pointer == 81 && y_pointer == 72)
||(x_pointer == 83 && y_pointer == 72)
||(x_pointer == 84 && y_pointer == 72)
||(x_pointer == 86 && y_pointer == 72)
||(x_pointer == 87 && y_pointer == 72)
||(x_pointer == 90 && y_pointer == 72)
||(x_pointer == 91 && y_pointer == 72)
||(x_pointer == 92 && y_pointer == 72)
||(x_pointer == 93 && y_pointer == 72)
||(x_pointer == 94 && y_pointer == 72)
||(x_pointer == 97 && y_pointer == 72)
||(x_pointer == 98 && y_pointer == 72)
||(x_pointer == 54 && y_pointer == 73)
||(x_pointer == 55 && y_pointer == 73)
||(x_pointer == 57 && y_pointer == 73)
||(x_pointer == 58 && y_pointer == 73)
||(x_pointer == 59 && y_pointer == 73)
||(x_pointer == 60 && y_pointer == 73)
||(x_pointer == 62 && y_pointer == 73)
||(x_pointer == 63 && y_pointer == 73)
||(x_pointer == 68 && y_pointer == 73)
||(x_pointer == 69 && y_pointer == 73)
||(x_pointer == 71 && y_pointer == 73)
||(x_pointer == 72 && y_pointer == 73)
||(x_pointer == 75 && y_pointer == 73)
||(x_pointer == 76 && y_pointer == 73)
||(x_pointer == 80 && y_pointer == 73)
||(x_pointer == 81 && y_pointer == 73)
||(x_pointer == 83 && y_pointer == 73)
||(x_pointer == 84 && y_pointer == 73)
||(x_pointer == 86 && y_pointer == 73)
||(x_pointer == 87 && y_pointer == 73)
||(x_pointer == 90 && y_pointer == 73)
||(x_pointer == 91 && y_pointer == 73)
||(x_pointer == 92 && y_pointer == 73)
||(x_pointer == 93 && y_pointer == 73)
||(x_pointer == 94 && y_pointer == 73)
||(x_pointer == 97 && y_pointer == 73)
||(x_pointer == 98 && y_pointer == 73)
||(x_pointer == 54 && y_pointer == 74)
||(x_pointer == 55 && y_pointer == 74)
||(x_pointer == 58 && y_pointer == 74)
||(x_pointer == 59 && y_pointer == 74)
||(x_pointer == 60 && y_pointer == 74)
||(x_pointer == 62 && y_pointer == 74)
||(x_pointer == 63 && y_pointer == 74)
||(x_pointer == 68 && y_pointer == 74)
||(x_pointer == 69 && y_pointer == 74)
||(x_pointer == 71 && y_pointer == 74)
||(x_pointer == 72 && y_pointer == 74)
||(x_pointer == 75 && y_pointer == 74)
||(x_pointer == 76 && y_pointer == 74)
||(x_pointer == 80 && y_pointer == 74)
||(x_pointer == 81 && y_pointer == 74)
||(x_pointer == 83 && y_pointer == 74)
||(x_pointer == 84 && y_pointer == 74)
||(x_pointer == 86 && y_pointer == 74)
||(x_pointer == 87 && y_pointer == 74)
||(x_pointer == 89 && y_pointer == 74)
||(x_pointer == 90 && y_pointer == 74)
||(x_pointer == 94 && y_pointer == 74)
||(x_pointer == 95 && y_pointer == 74)
||(x_pointer == 97 && y_pointer == 74)
||(x_pointer == 98 && y_pointer == 74)
||(x_pointer == 54 && y_pointer == 75)
||(x_pointer == 55 && y_pointer == 75)
||(x_pointer == 58 && y_pointer == 75)
||(x_pointer == 59 && y_pointer == 75)
||(x_pointer == 60 && y_pointer == 75)
||(x_pointer == 62 && y_pointer == 75)
||(x_pointer == 63 && y_pointer == 75)
||(x_pointer == 68 && y_pointer == 75)
||(x_pointer == 69 && y_pointer == 75)
||(x_pointer == 71 && y_pointer == 75)
||(x_pointer == 72 && y_pointer == 75)
||(x_pointer == 76 && y_pointer == 75)
||(x_pointer == 77 && y_pointer == 75)
||(x_pointer == 80 && y_pointer == 75)
||(x_pointer == 81 && y_pointer == 75)
||(x_pointer == 86 && y_pointer == 75)
||(x_pointer == 87 && y_pointer == 75)
||(x_pointer == 89 && y_pointer == 75)
||(x_pointer == 90 && y_pointer == 75)
||(x_pointer == 94 && y_pointer == 75)
||(x_pointer == 95 && y_pointer == 75)
||(x_pointer == 97 && y_pointer == 75)
||(x_pointer == 98 && y_pointer == 75)
||(x_pointer == 54 && y_pointer == 76)
||(x_pointer == 55 && y_pointer == 76)
||(x_pointer == 59 && y_pointer == 76)
||(x_pointer == 60 && y_pointer == 76)
||(x_pointer == 62 && y_pointer == 76)
||(x_pointer == 63 && y_pointer == 76)
||(x_pointer == 64 && y_pointer == 76)
||(x_pointer == 65 && y_pointer == 76)
||(x_pointer == 66 && y_pointer == 76)
||(x_pointer == 67 && y_pointer == 76)
||(x_pointer == 68 && y_pointer == 76)
||(x_pointer == 69 && y_pointer == 76)
||(x_pointer == 71 && y_pointer == 76)
||(x_pointer == 72 && y_pointer == 76)
||(x_pointer == 76 && y_pointer == 76)
||(x_pointer == 77 && y_pointer == 76)
||(x_pointer == 80 && y_pointer == 76)
||(x_pointer == 81 && y_pointer == 76)
||(x_pointer == 86 && y_pointer == 76)
||(x_pointer == 87 && y_pointer == 76)
||(x_pointer == 89 && y_pointer == 76)
||(x_pointer == 90 && y_pointer == 76)
||(x_pointer == 94 && y_pointer == 76)
||(x_pointer == 95 && y_pointer == 76)
||(x_pointer == 97 && y_pointer == 76)
||(x_pointer == 98 && y_pointer == 76)
||(x_pointer == 99 && y_pointer == 76)
||(x_pointer == 100 && y_pointer == 76)
||(x_pointer == 101 && y_pointer == 76)
||(x_pointer == 102 && y_pointer == 76))) || (main_difficulty == 4'd1 && ((x_pointer == 62 && y_pointer == 65)
||(x_pointer == 63 && y_pointer == 65)
||(x_pointer == 67 && y_pointer == 65)
||(x_pointer == 68 && y_pointer == 65)
||(x_pointer == 72 && y_pointer == 65)
||(x_pointer == 73 && y_pointer == 65)
||(x_pointer == 74 && y_pointer == 65)
||(x_pointer == 78 && y_pointer == 65)
||(x_pointer == 79 && y_pointer == 65)
||(x_pointer == 80 && y_pointer == 65)
||(x_pointer == 81 && y_pointer == 65)
||(x_pointer == 82 && y_pointer == 65)
||(x_pointer == 83 && y_pointer == 65)
||(x_pointer == 86 && y_pointer == 65)
||(x_pointer == 87 && y_pointer == 65)
||(x_pointer == 88 && y_pointer == 65)
||(x_pointer == 89 && y_pointer == 65)
||(x_pointer == 90 && y_pointer == 65)
||(x_pointer == 91 && y_pointer == 65)
||(x_pointer == 62 && y_pointer == 66)
||(x_pointer == 63 && y_pointer == 66)
||(x_pointer == 67 && y_pointer == 66)
||(x_pointer == 68 && y_pointer == 66)
||(x_pointer == 72 && y_pointer == 66)
||(x_pointer == 73 && y_pointer == 66)
||(x_pointer == 74 && y_pointer == 66)
||(x_pointer == 78 && y_pointer == 66)
||(x_pointer == 79 && y_pointer == 66)
||(x_pointer == 83 && y_pointer == 66)
||(x_pointer == 84 && y_pointer == 66)
||(x_pointer == 86 && y_pointer == 66)
||(x_pointer == 87 && y_pointer == 66)
||(x_pointer == 90 && y_pointer == 66)
||(x_pointer == 91 && y_pointer == 66)
||(x_pointer == 92 && y_pointer == 66)
||(x_pointer == 62 && y_pointer == 67)
||(x_pointer == 63 && y_pointer == 67)
||(x_pointer == 67 && y_pointer == 67)
||(x_pointer == 68 && y_pointer == 67)
||(x_pointer == 72 && y_pointer == 67)
||(x_pointer == 73 && y_pointer == 67)
||(x_pointer == 74 && y_pointer == 67)
||(x_pointer == 78 && y_pointer == 67)
||(x_pointer == 79 && y_pointer == 67)
||(x_pointer == 83 && y_pointer == 67)
||(x_pointer == 84 && y_pointer == 67)
||(x_pointer == 86 && y_pointer == 67)
||(x_pointer == 87 && y_pointer == 67)
||(x_pointer == 91 && y_pointer == 67)
||(x_pointer == 92 && y_pointer == 67)
||(x_pointer == 62 && y_pointer == 68)
||(x_pointer == 63 && y_pointer == 68)
||(x_pointer == 67 && y_pointer == 68)
||(x_pointer == 68 && y_pointer == 68)
||(x_pointer == 72 && y_pointer == 68)
||(x_pointer == 74 && y_pointer == 68)
||(x_pointer == 78 && y_pointer == 68)
||(x_pointer == 79 && y_pointer == 68)
||(x_pointer == 83 && y_pointer == 68)
||(x_pointer == 84 && y_pointer == 68)
||(x_pointer == 86 && y_pointer == 68)
||(x_pointer == 87 && y_pointer == 68)
||(x_pointer == 91 && y_pointer == 68)
||(x_pointer == 92 && y_pointer == 68)
||(x_pointer == 62 && y_pointer == 69)
||(x_pointer == 63 && y_pointer == 69)
||(x_pointer == 67 && y_pointer == 69)
||(x_pointer == 68 && y_pointer == 69)
||(x_pointer == 72 && y_pointer == 69)
||(x_pointer == 74 && y_pointer == 69)
||(x_pointer == 78 && y_pointer == 69)
||(x_pointer == 79 && y_pointer == 69)
||(x_pointer == 83 && y_pointer == 69)
||(x_pointer == 84 && y_pointer == 69)
||(x_pointer == 86 && y_pointer == 69)
||(x_pointer == 87 && y_pointer == 69)
||(x_pointer == 91 && y_pointer == 69)
||(x_pointer == 92 && y_pointer == 69)
||(x_pointer == 62 && y_pointer == 70)
||(x_pointer == 63 && y_pointer == 70)
||(x_pointer == 64 && y_pointer == 70)
||(x_pointer == 65 && y_pointer == 70)
||(x_pointer == 66 && y_pointer == 70)
||(x_pointer == 67 && y_pointer == 70)
||(x_pointer == 68 && y_pointer == 70)
||(x_pointer == 71 && y_pointer == 70)
||(x_pointer == 72 && y_pointer == 70)
||(x_pointer == 74 && y_pointer == 70)
||(x_pointer == 75 && y_pointer == 70)
||(x_pointer == 78 && y_pointer == 70)
||(x_pointer == 79 && y_pointer == 70)
||(x_pointer == 80 && y_pointer == 70)
||(x_pointer == 81 && y_pointer == 70)
||(x_pointer == 82 && y_pointer == 70)
||(x_pointer == 83 && y_pointer == 70)
||(x_pointer == 86 && y_pointer == 70)
||(x_pointer == 87 && y_pointer == 70)
||(x_pointer == 91 && y_pointer == 70)
||(x_pointer == 92 && y_pointer == 70)
||(x_pointer == 62 && y_pointer == 71)
||(x_pointer == 63 && y_pointer == 71)
||(x_pointer == 67 && y_pointer == 71)
||(x_pointer == 68 && y_pointer == 71)
||(x_pointer == 71 && y_pointer == 71)
||(x_pointer == 72 && y_pointer == 71)
||(x_pointer == 74 && y_pointer == 71)
||(x_pointer == 75 && y_pointer == 71)
||(x_pointer == 78 && y_pointer == 71)
||(x_pointer == 79 && y_pointer == 71)
||(x_pointer == 80 && y_pointer == 71)
||(x_pointer == 81 && y_pointer == 71)
||(x_pointer == 82 && y_pointer == 71)
||(x_pointer == 86 && y_pointer == 71)
||(x_pointer == 87 && y_pointer == 71)
||(x_pointer == 91 && y_pointer == 71)
||(x_pointer == 92 && y_pointer == 71)
||(x_pointer == 62 && y_pointer == 72)
||(x_pointer == 63 && y_pointer == 72)
||(x_pointer == 67 && y_pointer == 72)
||(x_pointer == 68 && y_pointer == 72)
||(x_pointer == 71 && y_pointer == 72)
||(x_pointer == 72 && y_pointer == 72)
||(x_pointer == 73 && y_pointer == 72)
||(x_pointer == 74 && y_pointer == 72)
||(x_pointer == 75 && y_pointer == 72)
||(x_pointer == 78 && y_pointer == 72)
||(x_pointer == 79 && y_pointer == 72)
||(x_pointer == 81 && y_pointer == 72)
||(x_pointer == 82 && y_pointer == 72)
||(x_pointer == 86 && y_pointer == 72)
||(x_pointer == 87 && y_pointer == 72)
||(x_pointer == 91 && y_pointer == 72)
||(x_pointer == 92 && y_pointer == 72)
||(x_pointer == 62 && y_pointer == 73)
||(x_pointer == 63 && y_pointer == 73)
||(x_pointer == 67 && y_pointer == 73)
||(x_pointer == 68 && y_pointer == 73)
||(x_pointer == 71 && y_pointer == 73)
||(x_pointer == 72 && y_pointer == 73)
||(x_pointer == 73 && y_pointer == 73)
||(x_pointer == 74 && y_pointer == 73)
||(x_pointer == 75 && y_pointer == 73)
||(x_pointer == 78 && y_pointer == 73)
||(x_pointer == 79 && y_pointer == 73)
||(x_pointer == 81 && y_pointer == 73)
||(x_pointer == 82 && y_pointer == 73)
||(x_pointer == 83 && y_pointer == 73)
||(x_pointer == 86 && y_pointer == 73)
||(x_pointer == 87 && y_pointer == 73)
||(x_pointer == 91 && y_pointer == 73)
||(x_pointer == 92 && y_pointer == 73)
||(x_pointer == 62 && y_pointer == 74)
||(x_pointer == 63 && y_pointer == 74)
||(x_pointer == 67 && y_pointer == 74)
||(x_pointer == 68 && y_pointer == 74)
||(x_pointer == 70 && y_pointer == 74)
||(x_pointer == 71 && y_pointer == 74)
||(x_pointer == 75 && y_pointer == 74)
||(x_pointer == 76 && y_pointer == 74)
||(x_pointer == 78 && y_pointer == 74)
||(x_pointer == 79 && y_pointer == 74)
||(x_pointer == 82 && y_pointer == 74)
||(x_pointer == 83 && y_pointer == 74)
||(x_pointer == 86 && y_pointer == 74)
||(x_pointer == 87 && y_pointer == 74)
||(x_pointer == 91 && y_pointer == 74)
||(x_pointer == 92 && y_pointer == 74)
||(x_pointer == 62 && y_pointer == 75)
||(x_pointer == 63 && y_pointer == 75)
||(x_pointer == 67 && y_pointer == 75)
||(x_pointer == 68 && y_pointer == 75)
||(x_pointer == 70 && y_pointer == 75)
||(x_pointer == 71 && y_pointer == 75)
||(x_pointer == 75 && y_pointer == 75)
||(x_pointer == 76 && y_pointer == 75)
||(x_pointer == 78 && y_pointer == 75)
||(x_pointer == 79 && y_pointer == 75)
||(x_pointer == 82 && y_pointer == 75)
||(x_pointer == 83 && y_pointer == 75)
||(x_pointer == 84 && y_pointer == 75)
||(x_pointer == 86 && y_pointer == 75)
||(x_pointer == 87 && y_pointer == 75)
||(x_pointer == 90 && y_pointer == 75)
||(x_pointer == 91 && y_pointer == 75)
||(x_pointer == 92 && y_pointer == 75)
||(x_pointer == 62 && y_pointer == 76)
||(x_pointer == 63 && y_pointer == 76)
||(x_pointer == 67 && y_pointer == 76)
||(x_pointer == 68 && y_pointer == 76)
||(x_pointer == 70 && y_pointer == 76)
||(x_pointer == 71 && y_pointer == 76)
||(x_pointer == 75 && y_pointer == 76)
||(x_pointer == 76 && y_pointer == 76)
||(x_pointer == 78 && y_pointer == 76)
||(x_pointer == 79 && y_pointer == 76)
||(x_pointer == 83 && y_pointer == 76)
||(x_pointer == 84 && y_pointer == 76)
||(x_pointer == 86 && y_pointer == 76)
||(x_pointer == 87 && y_pointer == 76)
||(x_pointer == 88 && y_pointer == 76)
||(x_pointer == 89 && y_pointer == 76)
||(x_pointer == 90 && y_pointer == 76)
||(x_pointer == 91 && y_pointer == 76)));
	wire level_display = (current_level == 0 && ((x_pointer == 94 && y_pointer == 41)
||(x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 99 && y_pointer == 41)
||(x_pointer == 100 && y_pointer == 41)
||(x_pointer == 94 && y_pointer == 42)
||(x_pointer == 95 && y_pointer == 42)
||(x_pointer == 99 && y_pointer == 42)
||(x_pointer == 100 && y_pointer == 42)
||(x_pointer == 94 && y_pointer == 43)
||(x_pointer == 95 && y_pointer == 43)
||(x_pointer == 99 && y_pointer == 43)
||(x_pointer == 100 && y_pointer == 43)
||(x_pointer == 94 && y_pointer == 44)
||(x_pointer == 95 && y_pointer == 44)
||(x_pointer == 99 && y_pointer == 44)
||(x_pointer == 100 && y_pointer == 44)
||(x_pointer == 94 && y_pointer == 45)
||(x_pointer == 95 && y_pointer == 45)
||(x_pointer == 99 && y_pointer == 45)
||(x_pointer == 100 && y_pointer == 45)
||(x_pointer == 94 && y_pointer == 46)
||(x_pointer == 95 && y_pointer == 46)
||(x_pointer == 99 && y_pointer == 46)
||(x_pointer == 100 && y_pointer == 46)
||(x_pointer == 94 && y_pointer == 47)
||(x_pointer == 95 && y_pointer == 47)
||(x_pointer == 99 && y_pointer == 47)
||(x_pointer == 100 && y_pointer == 47)
||(x_pointer == 94 && y_pointer == 48)
||(x_pointer == 95 && y_pointer == 48)
||(x_pointer == 99 && y_pointer == 48)
||(x_pointer == 100 && y_pointer == 48)
||(x_pointer == 94 && y_pointer == 49)
||(x_pointer == 95 && y_pointer == 49)
||(x_pointer == 99 && y_pointer == 49)
||(x_pointer == 100 && y_pointer == 49)
||(x_pointer == 94 && y_pointer == 50)
||(x_pointer == 95 && y_pointer == 50)
||(x_pointer == 99 && y_pointer == 50)
||(x_pointer == 100 && y_pointer == 50)
||(x_pointer == 94 && y_pointer == 51)
||(x_pointer == 95 && y_pointer == 51)
||(x_pointer == 96 && y_pointer == 51)
||(x_pointer == 97 && y_pointer == 51)
||(x_pointer == 98 && y_pointer == 51)
||(x_pointer == 99 && y_pointer == 51)
||(x_pointer == 100 && y_pointer == 51))) || (current_level == 1 && ((x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 42)
||(x_pointer == 97 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 96 && y_pointer == 43)
||(x_pointer == 97 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 97 && y_pointer == 44)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 97 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 97 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 97 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 97 && y_pointer == 49)
||(x_pointer == 98 && y_pointer == 49)
||(x_pointer == 97 && y_pointer == 50)
||(x_pointer == 98 && y_pointer == 50)
||(x_pointer == 97 && y_pointer == 51)
||(x_pointer == 98 && y_pointer == 51))) || (current_level == 2 && ((x_pointer == 94 && y_pointer == 41)
||(x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 99 && y_pointer == 41)
||(x_pointer == 94 && y_pointer == 42)
||(x_pointer == 95 && y_pointer == 42)
||(x_pointer == 96 && y_pointer == 42)
||(x_pointer == 97 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 99 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 99 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 99 && y_pointer == 44)
||(x_pointer == 94 && y_pointer == 45)
||(x_pointer == 95 && y_pointer == 45)
||(x_pointer == 96 && y_pointer == 45)
||(x_pointer == 97 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 99 && y_pointer == 45)
||(x_pointer == 94 && y_pointer == 46)
||(x_pointer == 95 && y_pointer == 46)
||(x_pointer == 96 && y_pointer == 46)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 99 && y_pointer == 46)
||(x_pointer == 94 && y_pointer == 47)
||(x_pointer == 95 && y_pointer == 47)
||(x_pointer == 94 && y_pointer == 48)
||(x_pointer == 95 && y_pointer == 48)
||(x_pointer == 94 && y_pointer == 49)
||(x_pointer == 95 && y_pointer == 49)
||(x_pointer == 94 && y_pointer == 50)
||(x_pointer == 95 && y_pointer == 50)
||(x_pointer == 96 && y_pointer == 50)
||(x_pointer == 97 && y_pointer == 50)
||(x_pointer == 98 && y_pointer == 50)
||(x_pointer == 99 && y_pointer == 50)
||(x_pointer == 94 && y_pointer == 51)
||(x_pointer == 95 && y_pointer == 51)
||(x_pointer == 96 && y_pointer == 51)
||(x_pointer == 97 && y_pointer == 51)
||(x_pointer == 98 && y_pointer == 51)
||(x_pointer == 99 && y_pointer == 51))) || (current_level == 3 && ((x_pointer == 94 && y_pointer == 41)
||(x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 99 && y_pointer == 41)
||(x_pointer == 94 && y_pointer == 42)
||(x_pointer == 95 && y_pointer == 42)
||(x_pointer == 96 && y_pointer == 42)
||(x_pointer == 97 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 99 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 99 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 99 && y_pointer == 44)
||(x_pointer == 94 && y_pointer == 45)
||(x_pointer == 95 && y_pointer == 45)
||(x_pointer == 96 && y_pointer == 45)
||(x_pointer == 97 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 99 && y_pointer == 45)
||(x_pointer == 94 && y_pointer == 46)
||(x_pointer == 95 && y_pointer == 46)
||(x_pointer == 96 && y_pointer == 46)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 99 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 99 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 99 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 49)
||(x_pointer == 99 && y_pointer == 49)
||(x_pointer == 94 && y_pointer == 50)
||(x_pointer == 95 && y_pointer == 50)
||(x_pointer == 96 && y_pointer == 50)
||(x_pointer == 97 && y_pointer == 50)
||(x_pointer == 98 && y_pointer == 50)
||(x_pointer == 99 && y_pointer == 50)
||(x_pointer == 94 && y_pointer == 51)
||(x_pointer == 95 && y_pointer == 51)
||(x_pointer == 96 && y_pointer == 51)
||(x_pointer == 97 && y_pointer == 51)
||(x_pointer == 98 && y_pointer == 51)
||(x_pointer == 99 && y_pointer == 51))) || (current_level == 4 && ((x_pointer == 97 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 42)
||(x_pointer == 96 && y_pointer == 43)
||(x_pointer == 96 && y_pointer == 44)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 95 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 95 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 94 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 94 && y_pointer == 48)
||(x_pointer == 95 && y_pointer == 48)
||(x_pointer == 96 && y_pointer == 48)
||(x_pointer == 97 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 99 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 49)
||(x_pointer == 98 && y_pointer == 50)
||(x_pointer == 98 && y_pointer == 51))) || (current_level == 5 && ((x_pointer == 94 && y_pointer == 41)
||(x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 94 && y_pointer == 42)
||(x_pointer == 94 && y_pointer == 43)
||(x_pointer == 94 && y_pointer == 44)
||(x_pointer == 94 && y_pointer == 45)
||(x_pointer == 94 && y_pointer == 46)
||(x_pointer == 95 && y_pointer == 46)
||(x_pointer == 96 && y_pointer == 46)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 49)
||(x_pointer == 94 && y_pointer == 50)
||(x_pointer == 98 && y_pointer == 50)
||(x_pointer == 95 && y_pointer == 51)
||(x_pointer == 96 && y_pointer == 51)
||(x_pointer == 97 && y_pointer == 51))) || (current_level == 6 && ((x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 94 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 94 && y_pointer == 43)
||(x_pointer == 94 && y_pointer == 44)
||(x_pointer == 94 && y_pointer == 45)
||(x_pointer == 95 && y_pointer == 45)
||(x_pointer == 96 && y_pointer == 45)
||(x_pointer == 97 && y_pointer == 45)
||(x_pointer == 94 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 94 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 94 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 94 && y_pointer == 49)
||(x_pointer == 98 && y_pointer == 49)
||(x_pointer == 94 && y_pointer == 50)
||(x_pointer == 98 && y_pointer == 50)
||(x_pointer == 95 && y_pointer == 51)
||(x_pointer == 96 && y_pointer == 51)
||(x_pointer == 97 && y_pointer == 51))) || (current_level == 7 && ((x_pointer == 94 && y_pointer == 41)
||(x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 99 && y_pointer == 41)
||(x_pointer == 94 && y_pointer == 42)
||(x_pointer == 95 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 99 && y_pointer == 42)
||(x_pointer == 94 && y_pointer == 43)
||(x_pointer == 95 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 99 && y_pointer == 43)
||(x_pointer == 97 && y_pointer == 44)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 99 && y_pointer == 44)
||(x_pointer == 97 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 96 && y_pointer == 47)
||(x_pointer == 97 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 96 && y_pointer == 48)
||(x_pointer == 97 && y_pointer == 48)
||(x_pointer == 96 && y_pointer == 49)
||(x_pointer == 97 && y_pointer == 49)
||(x_pointer == 96 && y_pointer == 50)
||(x_pointer == 97 && y_pointer == 50)
||(x_pointer == 95 && y_pointer == 51)
||(x_pointer == 96 && y_pointer == 51)
||(x_pointer == 97 && y_pointer == 51))) || (current_level == 8 && ((x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 94 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 94 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 94 && y_pointer == 44)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 94 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 95 && y_pointer == 46)
||(x_pointer == 96 && y_pointer == 46)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 94 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 94 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 94 && y_pointer == 49)
||(x_pointer == 98 && y_pointer == 49)
||(x_pointer == 94 && y_pointer == 50)
||(x_pointer == 98 && y_pointer == 50)
||(x_pointer == 95 && y_pointer == 51)
||(x_pointer == 96 && y_pointer == 51)
||(x_pointer == 97 && y_pointer == 51))) || (current_level == 9 && ((x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 94 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 94 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 94 && y_pointer == 44)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 94 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 94 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 95 && y_pointer == 47)
||(x_pointer == 96 && y_pointer == 47)
||(x_pointer == 97 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 49)
||(x_pointer == 94 && y_pointer == 50)
||(x_pointer == 98 && y_pointer == 50)
||(x_pointer == 95 && y_pointer == 51)
||(x_pointer == 96 && y_pointer == 51)
||(x_pointer == 97 && y_pointer == 51)));
endmodule